`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:52:26 03/31/2016 
// Design Name: 
// Module Name:    Deco_binaBCD 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Deco_binaBCD(
	input [6:0] Wr_bin,
	input sel_hora,SF_24_12,SF_AM_PM,
	output reg [7:0] Wr_BCD
    );

reg [7:0] Wr_BCD1;

always @*
	case (Wr_bin)
		7'b0000000: Wr_BCD1 = 8'b00000000;//00
		7'b0000001: Wr_BCD1 = 8'b00000001;//01
		7'b0000010: Wr_BCD1 = 8'b00000010;//02
		7'b0000011: Wr_BCD1 = 8'b00000011;//03
		7'b0000100: Wr_BCD1 = 8'b00000100;//04
		7'b0000101: Wr_BCD1 = 8'b00000101;//05
		7'b0000110: Wr_BCD1 = 8'b00000110;//06
		7'b0000111: Wr_BCD1 = 8'b00000111;//07
		7'b0001000: Wr_BCD1 = 8'b00001000;//08
		7'b0001001: Wr_BCD1 = 8'b00001001;//09
		7'b0001010: Wr_BCD1 = 8'b00010000;//10
		7'b0001011: Wr_BCD1 = 8'b00010001;//11
		7'b0001100: Wr_BCD1 = 8'b00010010;//12
		7'b0001101: Wr_BCD1 = 8'b00010011;//13
		7'b0001110: Wr_BCD1 = 8'b00010100;//14
		7'b0001111: Wr_BCD1 = 8'b00010101;//15
		7'b0010000: Wr_BCD1 = 8'b00010110;//16
		7'b0010001: Wr_BCD1 = 8'b00010111;//17
		7'b0010010: Wr_BCD1 = 8'b00011000;//18
		7'b0010011: Wr_BCD1 = 8'b00011001;//19
		7'b0010100: Wr_BCD1 = 8'b00100000;//20
		7'b0010101: Wr_BCD1 = 8'b00100001;//21
		7'b0010110: Wr_BCD1 = 8'b00100010;//22
		7'b0010111: Wr_BCD1 = 8'b00100011;//23
		7'b0011000: Wr_BCD1 = 8'b00100100;//24
		7'b0011001: Wr_BCD1 = 8'b00100101;//25
		7'b0011010: Wr_BCD1 = 8'b00100110;//26
		7'b0011011: Wr_BCD1 = 8'b00100111;//27
		7'b0011100: Wr_BCD1 = 8'b00101000;//28
		7'b0011101: Wr_BCD1 = 8'b00101001;//29
		7'b0011110: Wr_BCD1 = 8'b00110000;//30
		7'b0011111: Wr_BCD1 = 8'b00110001;//31
		7'b0100000: Wr_BCD1 = 8'b00110010;//32
		7'b0100001: Wr_BCD1 = 8'b00110011;//33
		7'b0100010: Wr_BCD1 = 8'b00110100;//34
		7'b0100011: Wr_BCD1 = 8'b00110101;//35
		7'b0100100: Wr_BCD1 = 8'b00110110;//36
		7'b0100101: Wr_BCD1 = 8'b00110111;//37
		7'b0100110: Wr_BCD1 = 8'b00111000;//38
		7'b0100111: Wr_BCD1 = 8'b00111001;//39
		7'b0101000: Wr_BCD1 = 8'b01000000;//40
		7'b0101001: Wr_BCD1 = 8'b01000001;//41
		7'b0101010: Wr_BCD1 = 8'b01000010;//42
		7'b0101011: Wr_BCD1 = 8'b01000011;//43
		7'b0101100: Wr_BCD1 = 8'b01000100;//44
		7'b0101101: Wr_BCD1 = 8'b01000101;//45
		7'b0101110: Wr_BCD1 = 8'b01000110;//46
		7'b0101111: Wr_BCD1 = 8'b01000111;//47
		7'b0110000: Wr_BCD1 = 8'b01001000;//48
		7'b0110001: Wr_BCD1 = 8'b01001001;//49
		7'b0110010: Wr_BCD1 = 8'b01010000;//50
		7'b0110011: Wr_BCD1 = 8'b01010001;//51
		7'b0110100: Wr_BCD1 = 8'b01010010;//52
		7'b0110101: Wr_BCD1 = 8'b01010011;//53
		7'b0110110: Wr_BCD1 = 8'b01010100;//54
		7'b0110111: Wr_BCD1 = 8'b01010101;//55
		7'b0111000: Wr_BCD1 = 8'b01010110;//56
		7'b0111001: Wr_BCD1 = 8'b01010111;//57
		7'b0111010: Wr_BCD1 = 8'b01011000;//58
		7'b0111011: Wr_BCD1 = 8'b01011001;//59
		7'b0111100: Wr_BCD1 = 8'b01100000;//60
		7'b0111101: Wr_BCD1 = 8'b01100001;//61
		7'b0111110: Wr_BCD1 = 8'b01100010;//62
		7'b0111111: Wr_BCD1 = 8'b01100011;//63
		7'b1000000: Wr_BCD1 = 8'b01100100;//64
		7'b1000001: Wr_BCD1 = 8'b01100101;//65
		7'b1000010: Wr_BCD1 = 8'b01100110;//66
		7'b1000011: Wr_BCD1 = 8'b01100111;//67
		7'b1000100: Wr_BCD1 = 8'b01101000;//68
		7'b1000101: Wr_BCD1 = 8'b01101001;//69
		7'b1000110: Wr_BCD1 = 8'b01110000;//70
		7'b1000111: Wr_BCD1 = 8'b01110001;//71
		7'b1001000: Wr_BCD1 = 8'b01110010;//72
		7'b1001001: Wr_BCD1 = 8'b01110011;//73
		7'b1001010: Wr_BCD1 = 8'b01110100;//74
		7'b1001011: Wr_BCD1 = 8'b01110101;//75
		7'b1001100: Wr_BCD1 = 8'b01110110;//76
		7'b1001101: Wr_BCD1 = 8'b01110111;//77
		7'b1001110: Wr_BCD1 = 8'b01111000;//78
		7'b1001111: Wr_BCD1 = 8'b01111001;//79
		7'b1010000: Wr_BCD1 = 8'b10000000;//80
		7'b1010001: Wr_BCD1 = 8'b10000001;//81
		7'b1010010: Wr_BCD1 = 8'b10000010;//82
		7'b1010011: Wr_BCD1 = 8'b10000011;//83
		7'b1010100: Wr_BCD1 = 8'b10000100;//84
		7'b1010101: Wr_BCD1 = 8'b10000101;//85
		7'b1010110: Wr_BCD1 = 8'b10000110;//86
		7'b1010111: Wr_BCD1 = 8'b10000111;//87
		7'b1011000: Wr_BCD1 = 8'b10001000;//88
		7'b1011001: Wr_BCD1 = 8'b10001001;//89
		7'b1011010: Wr_BCD1 = 8'b10010000;//90
		7'b1011011: Wr_BCD1 = 8'b10010001;//91
		7'b1011100: Wr_BCD1 = 8'b10010010;//92
		7'b1011101: Wr_BCD1 = 8'b10010011;//93
		7'b1011110: Wr_BCD1 = 8'b10010100;//94
		7'b1011111: Wr_BCD1 = 8'b10010101;//95
		7'b1100000: Wr_BCD1 = 8'b10010110;//96
		7'b1100001: Wr_BCD1 = 8'b10010111;//97
		7'b1100010: Wr_BCD1 = 8'b10011000;//98
		7'b1100011: Wr_BCD1 = 8'b10011001;//99
		7'b1100100: Wr_BCD1 = 8'b00000000;//00
		7'b1100101: Wr_BCD1 = 8'b00000000;//00
		7'b1100110: Wr_BCD1 = 8'b00000000;//00
		7'b1100111: Wr_BCD1 = 8'b00000000;//00
		7'b1101000: Wr_BCD1 = 8'b00000000;//00
		7'b1101001: Wr_BCD1 = 8'b00000000;//00
		7'b1101010: Wr_BCD1 = 8'b00000000;//00
		7'b1101011: Wr_BCD1 = 8'b00000000;//00
		7'b1101100: Wr_BCD1 = 8'b00000000;//00
		7'b1101101: Wr_BCD1 = 8'b00000000;//00
		7'b1101110: Wr_BCD1 = 8'b00000000;//00
		7'b1101111: Wr_BCD1 = 8'b00000000;//00
		7'b1110000: Wr_BCD1 = 8'b00000000;//00
		7'b1110001: Wr_BCD1 = 8'b00000000;//00
		7'b1110010: Wr_BCD1 = 8'b00000000;//00
		7'b1110011: Wr_BCD1 = 8'b00000000;//00
		7'b1110100: Wr_BCD1 = 8'b00000000;//00
		7'b1110101: Wr_BCD1 = 8'b00000000;//00
		7'b1110110: Wr_BCD1 = 8'b00000000;//00
		7'b1110111: Wr_BCD1 = 8'b00000000;//00
		7'b1111000: Wr_BCD1 = 8'b00000000;//00
		7'b1111001: Wr_BCD1 = 8'b00000000;//00
		7'b1111010: Wr_BCD1 = 8'b00000000;//00
		7'b1111011: Wr_BCD1 = 8'b00000000;//00
		7'b1111100: Wr_BCD1 = 8'b00000000;//00
		7'b1111101: Wr_BCD1 = 8'b00000000;//00
		7'b1111110: Wr_BCD1 = 8'b00000000;//00
		7'b1111111: Wr_BCD1 = 8'b00000000;//00
		default : Wr_BCD1 = 8'b00000000;//00
	endcase

always @*
	case ({sel_hora,SF_24_12})
		2'b00: Wr_BCD = Wr_BCD1;
		2'b01: Wr_BCD = Wr_BCD1;
		2'b10: Wr_BCD = Wr_BCD1;
		2'b11: Wr_BCD = {SF_AM_PM,Wr_BCD1[6:0]};
		default: Wr_BCD = Wr_BCD1;
	endcase
	
endmodule
